module data_memory(
    input [31:0] A,
    input [31:0] WD,
    input clk,
    input WE,
    output [31:0] RD
);

endmodule