module register_file(
    input [4:0] A1,
    input [4:0] A2,
    input [4:0] A3,
    input [31:0] WD3,
    input clk,
    input WE3,
    output [31:0] RD1,
    output [31:0] RD2
);
endmodule