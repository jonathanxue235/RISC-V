module instruction_memory(
    input [31:0] A,
    output [31:0] RD
);
    
   
endmodule